module score (
    input rst,
    input inGame,
    input hit,
    output reg [6:0] total;    
);

// 分出十位與個位給2個8*8 dot matrix 去顯示

endmodule //score