module DotMatrix (
    input clk_1khz,
    input rst,
    output reg [7:0] dot_col,
    output reg [7:0] dot_row
); // display total score

endmodule //DotMatrix